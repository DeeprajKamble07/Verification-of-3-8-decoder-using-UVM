interface intf;
  logic [2:0] a;
  logic [7:0] y;
endinterface
